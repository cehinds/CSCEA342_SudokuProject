`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: UAA Digital Circuits A342
// Engineer: Gwendolyn Beecher
// 
// Create Date: 11/30/2025 04:56:51 PM
// Design Name: VGA Sudoku Game
// Module Name: sudoku games
// Project Name: VGA Sudoku
//////////////////////////////////////////////////////////////////////////////////


module sudoku_puzzles(
    input  logic [1:0] selector,

    output logic [3:0] init_grid [0:8][0:8],
    output logic [3:0] solution  [0:8][0:8]
);

    logic [3:0] init_tmp [0:8][0:8];
    logic [3:0] sol_tmp  [0:8][0:8];

    // PUZZLE 1
    localparam logic [3:0] INIT1 [0:8][0:8] = '{
        '{5,3,0,0,7,0,0,0,0},
        '{6,0,0,1,9,5,0,0,0},
        '{0,9,8,0,0,0,0,6,0},
        '{8,0,0,0,6,0,0,0,3},
        '{4,0,0,8,0,3,0,0,1},
        '{7,0,0,0,2,0,0,0,6},
        '{0,6,0,0,0,0,2,8,0},
        '{0,0,0,4,1,9,0,0,5},
        '{0,0,0,0,8,0,0,7,9}
    };

    localparam logic [3:0] SOL1 [0:8][0:8] = '{
        '{5,3,4,6,7,8,9,1,2},
        '{6,7,2,1,9,5,3,4,8},
        '{1,9,8,3,4,2,5,6,7},
        '{8,5,9,7,6,1,4,2,3},
        '{4,2,6,8,5,3,7,9,1},
        '{7,1,3,9,2,4,8,5,6},
        '{9,6,1,5,3,7,2,8,4},
        '{2,8,7,4,1,9,6,3,5},
        '{3,4,5,2,8,6,1,7,9}
    };

    // PUZZLE 2
    localparam logic [3:0] INIT2 [0:8][0:8] = '{
        '{1,2,3,4,5,6,7,8,0},
        '{4,5,6,7,8,9,1,2,3},
        '{7,8,9,1,2,3,4,5,6},
        '{2,3,1,5,6,4,8,9,7},
        '{5,6,4,8,9,7,2,3,1},
        '{8,9,7,2,3,1,5,6,4},
        '{3,1,2,6,4,5,9,7,8},
        '{6,4,5,9,7,8,3,1,2},
        '{9,7,8,3,1,2,6,4,5}
    };

    localparam logic [3:0] SOL2 [0:8][0:8] = '{
        '{1,2,3,4,5,6,7,8,9},
        '{4,5,6,7,8,9,1,2,3},
        '{7,8,9,1,2,3,4,5,6},
        '{2,3,1,5,6,4,8,9,7},
        '{5,6,4,8,9,7,2,3,1},
        '{8,9,7,2,3,1,5,6,4},
        '{3,1,2,6,4,5,9,7,8},
        '{6,4,5,9,7,8,3,1,2},
        '{9,7,8,3,1,2,6,4,5}
    };

    // PUZZLE 3
    localparam logic [3:0] INIT3 [0:8][0:8] = '{
        '{0,0,0,2,6,0,7,0,1},
        '{6,8,0,0,7,0,0,9,0},
        '{1,9,0,0,0,4,5,0,0},
        '{8,2,0,1,0,0,0,4,0},
        '{0,4,0,6,0,2,9,0,0},
        '{0,5,0,0,0,3,0,2,8},
        '{0,9,0,3,0,0,0,7,4},
        '{0,4,0,0,5,0,0,3,6},
        '{7,0,3,0,1,8,0,0,0}
    };

    localparam logic [3:0] SOL3 [0:8][0:8] = '{
        '{4,3,5,2,6,9,7,8,1},
        '{6,8,2,5,7,1,4,9,3},
        '{1,9,7,8,3,4,5,6,2},
        '{8,2,6,1,9,5,3,4,7},
        '{3,7,4,6,8,2,9,1,5},
        '{9,5,1,7,4,3,6,2,8},
        '{5,1,9,3,2,6,8,7,4},
        '{2,4,8,9,5,7,1,3,6},
        '{7,6,3,4,1,8,2,5,9}
    };

    // Select puzzle
    always_comb begin
        case(selector)
            2'd0: begin init_tmp = INIT1; sol_tmp = SOL1; end
            2'd1: begin init_tmp = INIT2; sol_tmp = SOL2; end
            2'd2: begin init_tmp = INIT3; sol_tmp = SOL3; end
            default: begin init_tmp = INIT1; sol_tmp = SOL1; end
        endcase

        for (int r = 0; r < 9; r++)
            for (int c = 0; c < 9; c++) begin
                init_grid[r][c] = init_tmp[r][c];
                solution[r][c]  = sol_tmp[r][c];
            end
    end

endmodule
